---------------------------------------------------------------------
-- File Name: bubblesort.vhd
-- Project Name: Bubble sort algorithm
-- Decription: Implementation of bubble sort algorithm in FPGA
-- -----------------------------------------------------------------  
-- Author: Ritesh
-- email: ritesh.belgudri@gmail.com
-- Revision:
--
-- (c) 2018 https://github.com/riteshbel
---------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bubblesort is
port();
end entity bubblesort;

architecture rtl of bubblesort is


begin


end architecture rtl;
-- eof
