-- top file
