-- topfile
